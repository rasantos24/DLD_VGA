`timescale 1ns / 1ps
module Signal(
	input hcount,
	input vcount,
	output vsync,
	output hsync
    );

endmodule
