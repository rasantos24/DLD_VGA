
entity Signal is
end Signal;

architecture Behavioral of Signal is

begin


end Behavioral;

